module cl_adder_tb(
	input wire clk, Cout,
  	input wire [31:0] s,
  	output reg C0,
  	output reg [31:0] a, b);

endmodule