module comb_logic(
	input wire [7:0] input_data_in,
	output reg [7:0] output_data_out
);

endmodule
