module comb_logic(
input [7:0] input_wire,
output reg [7:0] output_wire);

endmodule
